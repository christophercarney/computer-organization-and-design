


module WBMux(

    );
endmodule
